module ReLu #(parameter )
(
    input clk,
    input activation_function,

);

  
      
