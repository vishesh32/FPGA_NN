`include "topology.sv"

module Neuron #(
    parameter

)

endmodule
